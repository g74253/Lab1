module ascii_decoder(
    input  logic [7:0] ascii_code,
    output logic [7:0] pattern [0:7]
);

    always_comb begin
        case (ascii_code)
            8'd65: // 'A'
                pattern = '{8'b00110000, 8'b01111000, 8'b11001100, 8'b11001100, 8'b11111100, 8'b11001100, 8'b11001100, 8'b00000000};
            8'd66: // 'B'
                pattern = '{8'b11111100, 8'b01100110, 8'b01100110, 8'b01111100, 8'b01100110, 8'b01100110, 8'b11111100, 8'b00000000};
            8'd67: // 'C'
                pattern = '{8'b00111100, 8'b01100110, 8'b11000000, 8'b11000000, 8'b11000000, 8'b01100110, 8'b00111100, 8'b00000000};
            8'd68: // 'D'
                pattern = '{8'b11111000, 8'b01101100, 8'b01100110, 8'b01100110, 8'b01100110, 8'b01101100, 8'b11111000, 8'b00000000};
            8'd69: // 'E'
                pattern = '{8'b11111110, 8'b01100010, 8'b01101000, 8'b01111000, 8'b01101000, 8'b01100010, 8'b11111110, 8'b00000000};
            8'd70: // 'F'
                pattern = '{8'b11111110, 8'b01100010, 8'b01101000, 8'b01111000, 8'b01101000, 8'b01100000, 8'b11110000, 8'b00000000};
            8'd71: // 'G'
                pattern = '{8'b00111100, 8'b01100110, 8'b11000000, 8'b11000000, 8'b11001110, 8'b01100110, 8'b00111110, 8'b00000000};
            8'd72: // 'H'
                pattern = '{8'b11001100, 8'b11001100, 8'b11001100, 8'b11111100, 8'b11001100, 8'b11001100, 8'b11001100, 8'b00000000};
            8'd73: // 'I'
                pattern = '{8'b01111000, 8'b00110000, 8'b00110000, 8'b00110000, 8'b00110000, 8'b00110000, 8'b01111000, 8'b00000000};
            8'd74: // 'J'
                pattern = '{8'b00011110, 8'b00001100, 8'b00001100, 8'b00001100, 8'b11001100, 8'b11001100, 8'b01111000, 8'b00000000};
            8'd75: // 'K'
                pattern = '{8'b11110110, 8'b01100110, 8'b01101100, 8'b01111000, 8'b01101100, 8'b01100110, 8'b11110110, 8'b00000000};
            8'd76: // 'L'
                pattern = '{8'b11110000, 8'b01100000, 8'b01100000, 8'b01100000, 8'b01100010, 8'b01100110, 8'b11111110, 8'b00000000};
            8'd77: // 'M'
                pattern = '{8'b11000110, 8'b11101110, 8'b11111110, 8'b11111110, 8'b11010110, 8'b11000110, 8'b11000110, 8'b00000000};
            8'd78: // 'N'
                pattern = '{8'b11000110, 8'b11100110, 8'b11110110, 8'b11011110, 8'b11001110, 8'b11000110, 8'b11000110, 8'b00000000};
            8'd79: // 'O'
                pattern = '{8'b00111000, 8'b01101100, 8'b11000110, 8'b11000110, 8'b11000110, 8'b01101100, 8'b00111000, 8'b00000000};
            8'd80: // 'P'
                pattern = '{8'b11111100, 8'b01100110, 8'b01100110, 8'b01111100, 8'b01100000, 8'b01100000, 8'b11110000, 8'b00000000};
            8'd81: // 'Q'
                pattern = '{8'b01111000, 8'b11001100, 8'b11001100, 8'b11001100, 8'b11011100, 8'b01111000, 8'b00011100, 8'b00000000};
            8'd82: // 'R'
                pattern = '{8'b11111100, 8'b01100110, 8'b01100110, 8'b01111100, 8'b01101100, 8'b01100110, 8'b11110110, 8'b00000000};
            8'd83: // 'S'
                pattern = '{8'b01111000, 8'b11001100, 8'b11100000, 8'b01110000, 8'b00011100, 8'b11001100, 8'b01111000, 8'b00000000};
            8'd84: // 'T'
                pattern = '{8'b11111100, 8'b10110100, 8'b00110000, 8'b00110000, 8'b00110000, 8'b00110000, 8'b01111000, 8'b00000000};
            8'd85: // 'U'
                pattern = '{8'b11001100, 8'b11001100, 8'b11001100, 8'b11001100, 8'b11001100, 8'b11001100, 8'b11111100, 8'b00000000};
            8'd86: // 'V'
                pattern = '{8'b11001100, 8'b11001100, 8'b11001100, 8'b11001100, 8'b11001100, 8'b01111000, 8'b00110000, 8'b00000000};
            8'd87: // 'W'
                pattern = '{8'b11000110, 8'b11000110, 8'b11000110, 8'b11010110, 8'b11111110, 8'b11101110, 8'b11000110, 8'b00000000};
            8'd88: // 'X'
                pattern = '{8'b11000110, 8'b11000110, 8'b01101100, 8'b00111000, 8'b00111000, 8'b01101100, 8'b11000110, 8'b00000000};
            8'd89: // 'Y'
                pattern = '{8'b11001100, 8'b11001100, 8'b11001100, 8'b01111000, 8'b00110000, 8'b00110000, 8'b01111000, 8'b00000000};
            8'd90: // 'Z'
                pattern = '{8'b11111110, 8'b11000110, 8'b10001100, 8'b00011000, 8'b00110010, 8'b01100110, 8'b11111110, 8'b00000000};
					 
				8'd48: // '0'
					 pattern = '{8'b01111000, 8'b11001100, 8'b11011100, 8'b11111100, 8'b11101100, 8'b11001100, 8'b01111100, 8'b00000000};
				8'd49: // '1'
					 pattern = '{8'b00110000, 8'b01110000, 8'b00110000, 8'b00110000, 8'b00110000, 8'b00110000, 8'b11111100, 8'b00000000};
				8'd50: // '2'
					 pattern = '{8'b01111000, 8'b11001100, 8'b00001100, 8'b00111000, 8'b01100000, 8'b11001100, 8'b11111100, 8'b00000000};
				8'd51: // '3'
					 pattern = '{8'b01111000, 8'b11001100, 8'b00001100, 8'b00111000, 8'b00001100, 8'b11001100, 8'b01111000, 8'b00000000};
				8'd52: // '4'
					 pattern = '{8'b00011100, 8'b00111100, 8'b01101100, 8'b11001100, 8'b11111110, 8'b00001100, 8'b00011110, 8'b00000000};
				8'd53: // '5'
					 pattern = '{8'b11111100, 8'b11000000, 8'b11111000, 8'b00001100, 8'b00001100, 8'b11001100, 8'b01111000, 8'b00000000};
				8'd54: // '6'
					 pattern = '{8'b00111000, 8'b01100000, 8'b11000000, 8'b11111000, 8'b11001100, 8'b11001100, 8'b01111000, 8'b00000000};
				8'd55: // '7'
					 pattern = '{8'b11111100, 8'b11001100, 8'b00001100, 8'b00011000, 8'b00110000, 8'b00110000, 8'b00110000, 8'b00000000};
				8'd56: // '8'
					 pattern = '{8'b01111000, 8'b11001100, 8'b11001100, 8'b01111000, 8'b11001100, 8'b11001100, 8'b01111000, 8'b00000000};
				8'd57: // '9'
					 pattern = '{8'b01111000, 8'b11001100, 8'b11001100, 8'b01111100, 8'b00001100, 8'b00011000, 8'b01110000, 8'b00000000};
					 

				8'd97: // 'a'
					 pattern = '{8'b00000000, 8'b00000000, 8'b01111000, 8'b00001100, 8'b01111100, 8'b11001100, 8'b01110110, 8'b00000000};
				8'd98: // 'b'
					 pattern = '{8'b11100000, 8'b01100000, 8'b01100000, 8'b01111100, 8'b01100110, 8'b01100110, 8'b11011100, 8'b00000000};
				8'd99: // 'c'
					 pattern = '{8'b00000000, 8'b00000000, 8'b01111000, 8'b11001100, 8'b11000000, 8'b11001100, 8'b01111000, 8'b00000000};
				8'd100: // 'd'
					 pattern = '{8'b00011100, 8'b00001100, 8'b00001100, 8'b01111100, 8'b11001100, 8'b11001100, 8'b01110110, 8'b00000000};
				8'd101: // 'e'
					 pattern = '{8'b00000000, 8'b00000000, 8'b01111000, 8'b11001100, 8'b11111100, 8'b11000000, 8'b01111000, 8'b00000000};
				8'd102: // 'f'
					 pattern = '{8'b00111000, 8'b01101100, 8'b01100000, 8'b11110000, 8'b01100000, 8'b01100000, 8'b11110000, 8'b00000000};
				8'd103: // 'g'
					 pattern = '{8'b00000000, 8'b00000000, 8'b01110110, 8'b11001100, 8'b11001100, 8'b01111100, 8'b00001100, 8'b11111000};
				8'd104: // 'h'
					 pattern = '{8'b11100000, 8'b01100000, 8'b01101100, 8'b01110110, 8'b01100110, 8'b01100110, 8'b11100110, 8'b00000000};
				8'd105: // 'i'
					 pattern = '{8'b00110000, 8'b00000000, 8'b01110000, 8'b00110000, 8'b00110000, 8'b00110000, 8'b01111000, 8'b00000000};
				8'd106: // 'j'
					 pattern = '{8'b00001100, 8'b00000000, 8'b00001100, 8'b00001100, 8'b00001100, 8'b11001100, 8'b11001100, 8'b01111000};
				8'd107: // 'k'
					 pattern = '{8'b11100000, 8'b01100000, 8'b01100110, 8'b01101100, 8'b01111000, 8'b01101100, 8'b11100110, 8'b00000000};
				8'd108: // 'l'
					 pattern = '{8'b01110000, 8'b00110000, 8'b00110000, 8'b00110000, 8'b00110000, 8'b00110000, 8'b01111000, 8'b00000000};
				8'd109: // 'm'
					 pattern = '{8'b00000000, 8'b00000000, 8'b11001100, 8'b11111110, 8'b11111110, 8'b11010110, 8'b11000110, 8'b00000000};
				8'd110: // 'n'
					 pattern = '{8'b00000000, 8'b00000000, 8'b11111000, 8'b11001100, 8'b11001100, 8'b11001100, 8'b11001100, 8'b00000000};
				8'd111: // 'o'
					 pattern = '{8'b00000000, 8'b00000000, 8'b01111000, 8'b11001100, 8'b11001100, 8'b11001100, 8'b01111000, 8'b00000000};
				8'd112: // 'p'
					 pattern = '{8'b00000000, 8'b00000000, 8'b11011100, 8'b01100110, 8'b01100110, 8'b01111100, 8'b01100000, 8'b11110000};
				8'd113: // 'q'
					 pattern = '{8'b00000000, 8'b00000000, 8'b01110110, 8'b11001100, 8'b11001100, 8'b01111100, 8'b00001100, 8'b00011110};
				8'd114: // 'r'
					 pattern = '{8'b00000000, 8'b00000000, 8'b10011100, 8'b01110110, 8'b01100110, 8'b01100000, 8'b11110000, 8'b00000000};
				8'd115: // 's'
					 pattern = '{8'b00000000, 8'b00000000, 8'b01111100, 8'b11000000, 8'b01111000, 8'b00001100, 8'b11111000, 8'b00000000};
				8'd116: // 't'
					 pattern = '{8'b00010000, 8'b00110000, 8'b01111100, 8'b00110000, 8'b00110000, 8'b00110100, 8'b00011000, 8'b00000000};
				8'd117: // 'u'
					 pattern = '{8'b00000000, 8'b00000000, 8'b11001100, 8'b11001100, 8'b11001100, 8'b11001100, 8'b01110110, 8'b00000000};
				8'd118: // 'v'
					 pattern = '{8'b00000000, 8'b00000000, 8'b11001100, 8'b11001100, 8'b11001100, 8'b01111000, 8'b00110000, 8'b00000000};
				8'd119: // 'w'
					 pattern = '{8'b00000000, 8'b00000000, 8'b11000110, 8'b11000110, 8'b11010110, 8'b11111110, 8'b01101100, 8'b00000000};
				8'd120: // 'x'
					 pattern = '{8'b00000000, 8'b00000000, 8'b11000110, 8'b01101100, 8'b00111000, 8'b01101100, 8'b11000110, 8'b00000000};
				8'd121: // 'y'
					 pattern = '{8'b00000000, 8'b00000000, 8'b11001100, 8'b11001100, 8'b11001100, 8'b01111100, 8'b00001100, 8'b11111000};
				8'd122: // 'z'
					 pattern = '{8'b00000000, 8'b00000000, 8'b11111100, 8'b10011000, 8'b00110000, 8'b01100100, 8'b11111100, 8'b00000000};

					 
					 
            default: // default case for unsupported characters
                pattern = '{default: 8'b00000000};
        endcase
    end

endmodule
