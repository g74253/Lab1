module decodificador(
    input [3:0] e,
    output [6:0] c
);

assign c = (e == 4'b0000) ? 7'b1000000 :
           (e == 4'b0001) ? 7'b1111001 :
           (e == 4'b0010) ? 7'b0100100 :
           (e == 4'b0011) ? 7'b0110000 :
           (e == 4'b0100) ? 7'b0011001 :
           (e == 4'b0101) ? 7'b0010010 :
           (e == 4'b0110) ? 7'b0000010 :
           (e == 4'b0111) ? 7'b1111000 :
           (e == 4'b1000) ? 7'b0000000 :
           (e == 4'b1001) ? 7'b0011000 :
           (e == 4'b1010) ? 7'b0001000 :
           (e == 4'b1011) ? 7'b0000011 :
           (e == 4'b1100) ? 7'b1000110 :
           (e == 4'b1101) ? 7'b0100001 :
           (e == 4'b1110) ? 7'b0000110 :
           (e == 4'b1111) ? 7'b0001110 :
                            7'b0100100;

endmodule