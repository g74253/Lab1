module setup(input logic end_setup
				input logic boton_arriba,
				input logic boton_abajo,
				input logic boton_izquierda,
				input logic boton_derecha,
				input logic [2:0] cant_barco,
				input logic matriz,
				input logic boton_colocar);
				
				
				
	always @()begin
	end
endmodule